*Current mirror

*.include 180nm.lib
*.include tsmc018p.lib
.MODEL  CMOSN NMOS LEVEL=1 KP=5E-005 VT0=.7 LAMBDA=0.01

.MODEL  CMOSP PMOS LEVEL=1 KP=2E-005 VT0=-.7 LAMBDA=0.01

M1 2 2 1 1 CMOSP l=1.2u w=9000n
M2 3 2 1 1 CMOSP l=1.2u w=9000n
M3 3 4 0 0 CMOSN l=1.2u w = {w}
C1 3 0 100p
ICM 2 0 500u
VDD 1 0 5
Vsig 4 5 ac sin(0 10m 1k)
Vdc 5 0 2
*.op
*.dc Vdc 0 5 0.05; DC level
.param w = 2u
.step param w 10u 14u 0.5u
.ac dec 10 1 1g
.end


