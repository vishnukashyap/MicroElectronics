**clipper circuit**

.model DIN4007 D (IS=7.02767e-09 RS=0.0341512 N=1.80803 EG=1.05743 XTI=5 BV=1000 IBV=5e-08 CJO=1e-11 VJ=0.7 M=0.5 FC=0.5 TT=1e-07 KF=0 AF=1)

V1 1 0 sin(0 5 1)
R1 1 2 1k
D1 0 2 DIN4007


*.op
.tran 1 10 0
.end

