VCVS

Rs 1 2 100
Ri 2 0 2Meg
Ro 3 4 100
Cl 4 0 100n

Vin 1 0 ac sin(1 50m 1k)
E1 3 0 2 0 100

*.op
*.tran 1m 10m
*.four 1k V(4) I(Ro) I(E1) I(Vin)
*.ac dec 10 1 100Meg

*.noise is used to find the noise signals introduced in the circuit by the electrical components. It's syntax is .noise followed by the output node at which you calculate the noise, the input source, analysis type (lin/oct/dec), number of points in each unit, starting frequency and stopping frequency.
.noise V(4) Vin dec 10 1 1Meg
