**current miror**
.MODEL CMOSN NMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 4.1E-9
+XJ      = 1E-7           NCH     = 2.3549E17      VTH0    = 0.3694303
+K1      = 0.5789116      K2      = 1.110723E-3    K3      = 1E-3
+K3B     = 0.0297124      W0      = 1E-7           NLX     = 2.037748E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 1.2953626      DVT1    = 0.3421545      DVT2    = 0.0395588
+U0      = 293.1687573    UA      = -1.21942E-9    UB      = 2.325738E-18
+UC      = 7.061289E-11   VSAT    = 1.676164E5     A0      = 2
+AGS     = 0.4764546      B0      = 1.617101E-7    B1      = 5E-6
+KETA    = -0.0138552     A1      = 1.09168E-3     A2      = 0.3303025
+RDSW    = 105.6133217    PRWG    = 0.5            PRWB    = -0.2
+WR      = 1              WINT    = 2.885735E-9    LINT    = 1.715622E-8
+XL      = 0              XW      = -1E-8          DWG     = 2.754317E-9
+DWB     = -3.690793E-9   VOFF    = -0.0948017     NFACTOR = 2.1860065
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 2.665034E-3    ETAB    = 6.028975E-5
+DSUB    = 0.0442223      PCLM    = 1.746064       PDIBLC1 = 0.3258185
+PDIBLC2 = 2.701992E-3    PDIBLCB = -0.1           DROUT   = 0.9787232
+PSCBE1  = 4.494778E10    PSCBE2  = 3.672074E-8    PVAG    = 0.0122755
+DELTA   = 0.01           RSH     = 7              MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 8.58E-10       CGSO    = 8.58E-10       CGBO    = 1E-12
+CJ      = 9.471097E-4    PB      = 0.8            MJ      = 0.3726161
+CJSW    = 1.905901E-10   PBSW    = 0.8            MJSW    = 0.1369758
+CJSWG   = 3.3E-10        PBSWG   = 0.8            MJSWG   = 0.1369758
+CF      = 0              PVTH0   = -5.105777E-3   PRDSW   = -1.1011726
+PK2     = 2.247806E-3    WKETA   = -5.071892E-3   LKETA   = 5.324922E-4
+PU0     = -4.0206081     PUA     = -4.48232E-11   PUB     = 5.018589E-24
+PVSAT   = 2E3            PETA0   = 1E-4           PKETA   = -2.090695E-3    )
*
.MODEL CMOSP PMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 4.1E-9
+XJ      = 1E-7           NCH     = 4.1589E17      VTH0    = -0.3823437
+K1      = 0.5722049      K2      = 0.0219717      K3      = 0.1576753
+K3B     = 4.2763642      W0      = 1E-6           NLX     = 1.104212E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 0.6234839      DVT1    = 0.2479255      DVT2    = 0.1
+U0      = 109.4682454    UA      = 1.31646E-9     UB      = 1E-21
+UC      = -1E-10         VSAT    = 1.054892E5     A0      = 1.5796859
+AGS     = 0.3115024      B0      = 4.729297E-7    B1      = 1.446715E-6
+KETA    = 0.0298609      A1      = 0.3886886      A2      = 0.4010376
+RDSW    = 199.1594405    PRWG    = 0.5            PRWB    = -0.4947034
+WR      = 1              WINT    = 0              LINT    = 2.93948E-8
+XL      = 0              XW      = -1E-8          DWG     = -1.998034E-8
+DWB     = -2.481453E-9   VOFF    = -0.0935653     NFACTOR = 2
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 3.515392E-4    ETAB    = -4.804338E-4
+DSUB    = 1.215087E-5    PCLM    = 0.96422        PDIBLC1 = 3.026627E-3
+PDIBLC2 = -1E-5          PDIBLCB = -1E-3          DROUT   = 1.117016E-4
+PSCBE1  = 7.999986E10    PSCBE2  = 8.271897E-10   PVAG    = 0.0190118
+DELTA   = 0.01           RSH     = 8.1            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 7.82E-10       CGSO    = 7.82E-10       CGBO    = 1E-12
+CJ      = 1.214428E-3    PB      = 0.8461606      MJ      = 0.4192076
+CJSW    = 2.165642E-10   PBSW    = 0.8            MJSW    = 0.3202874
+CJSWG   = 4.22E-10       PBSWG   = 0.8            MJSWG   = 0.3202874
+CF      = 0              PVTH0   = 5.167913E-4    PRDSW   = 9.5068821
+PK2     = 1.095907E-3    WKETA   = 0.0133232      LKETA   = -3.648003E-3
+PU0     = -1.0674346     PUA     = -4.30826E-11   PUB     = 1E-21
+PVSAT   = 50             PETA0   = 1E-4           PKETA   = -1.822724E-3    )
*
Vdd 4 0 3.3
Iref 2 1 10u
M1 1 1 0 0 CMOSN L=10u W=10u
M2 3 1 0 0 CMOSN L=10u W=100u
V1 3 0 3.3
R1 4 2 {R}
*R1 4 2 100k
*.op
.step param R 100k 500k 50k
.dc V1 0 3.3 0.1
